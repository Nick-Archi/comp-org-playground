module myControlUnit();

endmodule